`timescale 1ns / 1ns
`include "Problem22.v"

module shift_register8_tb;

	reg [7:0] Din;
	reg clk;
	wire [7:0] Qout

endmodule
