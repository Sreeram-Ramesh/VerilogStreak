// Modelling a Inverter

module top_module (in_1, out_1);

    input in_1;
    output out_1;

    assign out_1 = ~in_1;

endmodule
